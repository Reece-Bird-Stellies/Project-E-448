*********************************************************************
//--- Inductors ---
L1     1   2  -
//----- Ports -----
P1     1   0
P2     2   0
.end
